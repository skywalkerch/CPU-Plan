library verilog;
use verilog.vl_types.all;
entity nandTest is
    port(
        Pop             : out    vl_logic;
        Pid             : out    vl_logic
    );
end nandTest;
