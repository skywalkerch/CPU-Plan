library verilog;
use verilog.vl_types.all;
entity nandTest_vlg_vec_tst is
end nandTest_vlg_vec_tst;
