library verilog;
use verilog.vl_types.all;
entity CLA4_vlg_vec_tst is
end CLA4_vlg_vec_tst;
